module main

import json112

fn main(){
	s := '{"name":"aaa"}'
	json112.decode(s)	
}