module json112

fn utf16str_to_unicodepoint(str string,pos int)?Unicode{
	return Unicode{}
}