module json112

[if jsondebug]
fn log<T>(msg T){
	println(msg)
}